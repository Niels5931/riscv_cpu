library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity riscv_cpu_tb is
end entity;

architecture tb of riscv_cpu_tb is

	begin

end architecture;
