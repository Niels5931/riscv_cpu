library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ins_mem_tb is
end entity;

architecture tb of ins_mem_tb is

	begin

end architecture;
