library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity package_tb is
end entity;

architecture tb of package_tb is

	begin

end architecture;
